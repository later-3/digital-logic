module adder (
 input a,b,
 output [1:0] sum
);
 assign sum=a+b;
endmodule
